magic
tech sky130A
timestamp 1743308394
<< nwell >>
rect -70 95 200 535
<< nmos >>
rect 50 -60 65 40
rect 115 -60 130 40
<< pmos >>
rect 50 115 65 515
rect 115 115 130 515
<< ndiff >>
rect 0 25 50 40
rect 0 -45 15 25
rect 35 -45 50 25
rect 0 -60 50 -45
rect 65 25 115 40
rect 65 -45 80 25
rect 100 -45 115 25
rect 65 -60 115 -45
rect 130 25 180 40
rect 130 -45 145 25
rect 165 -45 180 25
rect 130 -60 180 -45
<< pdiff >>
rect 0 500 50 515
rect 0 130 15 500
rect 35 130 50 500
rect 0 115 50 130
rect 65 115 115 515
rect 130 500 180 515
rect 130 130 145 500
rect 165 130 180 500
rect 130 115 180 130
<< ndiffc >>
rect 15 -45 35 25
rect 80 -45 100 25
rect 145 -45 165 25
<< pdiffc >>
rect 15 130 35 500
rect 145 130 165 500
<< psubdiff >>
rect -50 25 0 40
rect -50 -45 -35 25
rect -15 -45 0 25
rect -50 -60 0 -45
<< nsubdiff >>
rect -50 500 0 515
rect -50 130 -35 500
rect -15 130 0 500
rect -50 115 0 130
<< psubdiffcont >>
rect -35 -45 -15 25
<< nsubdiffcont >>
rect -35 130 -15 500
<< poly >>
rect 50 515 65 530
rect 115 515 130 530
rect 50 95 65 115
rect 10 85 65 95
rect 10 65 20 85
rect 40 65 65 85
rect 10 55 65 65
rect 50 40 65 55
rect 115 95 130 115
rect 115 85 170 95
rect 115 65 140 85
rect 160 65 170 85
rect 115 55 170 65
rect 115 40 130 55
rect 50 -75 65 -60
rect 115 -75 130 -60
<< polycont >>
rect 20 65 40 85
rect 140 65 160 85
<< locali >>
rect -45 565 45 575
rect -45 545 -35 565
rect -15 545 15 565
rect 35 545 45 565
rect -45 500 45 545
rect -45 130 -35 500
rect -15 130 15 500
rect 35 130 45 500
rect 135 500 175 510
rect 135 160 145 500
rect -45 120 45 130
rect 70 130 145 160
rect 165 130 175 500
rect 70 120 175 130
rect 10 85 50 95
rect 10 65 20 85
rect 40 65 50 85
rect 10 55 50 65
rect 70 85 110 120
rect 70 65 80 85
rect 100 65 110 85
rect -45 25 45 35
rect -45 -45 -35 25
rect -15 -45 15 25
rect 35 -45 45 25
rect -45 -90 45 -45
rect 70 25 110 65
rect 130 85 170 95
rect 130 65 140 85
rect 160 65 170 85
rect 130 55 170 65
rect 70 -45 80 25
rect 100 -45 110 25
rect 70 -55 110 -45
rect 135 25 175 35
rect 135 -45 145 25
rect 165 -45 175 25
rect -45 -110 -35 -90
rect -15 -110 15 -90
rect 35 -110 45 -90
rect -45 -120 45 -110
rect 135 -90 175 -45
rect 135 -110 145 -90
rect 165 -110 175 -90
rect 135 -120 175 -110
<< viali >>
rect -35 545 -15 565
rect 15 545 35 565
rect 20 65 40 85
rect 80 65 100 85
rect 140 65 160 85
rect -35 -110 -15 -90
rect 15 -110 35 -90
rect 145 -110 165 -90
<< metal1 >>
rect -70 565 200 575
rect -70 545 -35 565
rect -15 545 15 565
rect 35 545 200 565
rect -70 535 200 545
rect 10 85 50 95
rect 10 65 20 85
rect 40 65 50 85
rect 10 55 50 65
rect 70 85 110 95
rect 70 65 80 85
rect 100 65 110 85
rect 70 55 110 65
rect 130 85 170 95
rect 130 65 140 85
rect 160 65 170 85
rect 130 55 170 65
rect -70 -90 200 -80
rect -70 -110 -35 -90
rect -15 -110 15 -90
rect 35 -110 145 -90
rect 165 -110 200 -90
rect -70 -120 200 -110
<< labels >>
flabel metal1 10 75 10 75 7 FreeSans 80 0 -40 0 A
port 1 w
flabel metal1 170 75 170 75 3 FreeSans 80 0 40 0 B
port 2 e
flabel metal1 70 75 70 75 7 FreeSans 80 0 -40 0 Y
port 3 w
flabel metal1 -70 -100 -70 -100 7 FreeSans 80 0 -40 0 GND
port 5 w
flabel metal1 -70 555 -70 555 7 FreeSans 80 0 -40 0 VDD
port 4 w
<< end >>
