magic
tech sky130A
timestamp 1743203493
<< nwell >>
rect -70 95 200 240
<< nmos >>
rect 50 -50 65 50
rect 115 -50 130 50
<< pmos >>
rect 50 115 65 215
rect 115 115 130 215
<< ndiff >>
rect 0 35 50 50
rect 0 -35 15 35
rect 35 -35 50 35
rect 0 -50 50 -35
rect 65 -50 115 50
rect 130 35 180 50
rect 130 -35 145 35
rect 165 -35 180 35
rect 130 -50 180 -35
<< pdiff >>
rect 0 200 50 215
rect 0 130 15 200
rect 35 130 50 200
rect 0 115 50 130
rect 65 200 115 215
rect 65 130 80 200
rect 100 130 115 200
rect 65 115 115 130
rect 130 200 180 215
rect 130 130 145 200
rect 165 130 180 200
rect 130 115 180 130
<< ndiffc >>
rect 15 -35 35 35
rect 145 -35 165 35
<< pdiffc >>
rect 15 130 35 200
rect 80 130 100 200
rect 145 130 165 200
<< psubdiff >>
rect -50 35 0 50
rect -50 -35 -35 35
rect -15 -35 0 35
rect -50 -50 0 -35
<< nsubdiff >>
rect -50 200 0 215
rect -50 130 -35 200
rect -15 130 0 200
rect -50 115 0 130
<< psubdiffcont >>
rect -35 -35 -15 35
<< nsubdiffcont >>
rect -35 130 -15 200
<< poly >>
rect 50 215 65 230
rect 115 215 130 230
rect 50 50 65 115
rect 115 50 130 115
rect 50 -65 65 -50
rect 115 -65 130 -50
rect 25 -75 65 -65
rect 25 -95 35 -75
rect 55 -95 65 -75
rect 25 -105 65 -95
rect 90 -75 130 -65
rect 90 -95 100 -75
rect 120 -95 130 -75
rect 90 -105 130 -95
<< polycont >>
rect 35 -95 55 -75
rect 100 -95 120 -75
<< locali >>
rect -45 200 45 210
rect -45 130 -35 200
rect -15 130 15 200
rect 35 130 45 200
rect -45 120 45 130
rect 70 200 110 210
rect 70 130 80 200
rect 100 130 110 200
rect 70 120 110 130
rect 135 200 175 210
rect 135 130 145 200
rect 165 130 175 200
rect 135 120 175 130
rect 90 90 110 120
rect 90 70 200 90
rect 155 45 175 70
rect -45 35 45 45
rect -45 -35 -35 35
rect -15 -35 15 35
rect 35 -35 45 35
rect -45 -45 45 -35
rect 135 35 175 45
rect 135 -35 145 35
rect 165 -35 175 35
rect 135 -45 175 -35
rect -70 -75 65 -65
rect -70 -85 35 -75
rect 25 -95 35 -85
rect 55 -95 65 -75
rect 25 -105 65 -95
rect 90 -75 130 -65
rect 90 -95 100 -75
rect 120 -95 130 -75
rect 90 -105 130 -95
rect 105 -125 130 -105
rect -70 -145 130 -125
<< viali >>
rect -35 130 -15 200
rect 15 130 35 200
rect 145 130 165 200
rect -35 -35 -15 35
rect 15 -35 35 35
<< metal1 >>
rect -70 200 200 210
rect -70 130 -35 200
rect -15 130 15 200
rect 35 130 145 200
rect 165 130 200 200
rect -70 120 200 130
rect -70 35 200 45
rect -70 -35 -35 35
rect -15 -35 15 35
rect 35 -35 200 35
rect -70 -45 200 -35
<< labels >>
flabel locali -70 -135 -70 -135 7 FreeSans 80 0 -40 0 B
port 2 w
flabel locali -70 -75 -70 -75 7 FreeSans 80 0 -40 0 A
port 1 w
flabel metal1 -70 0 -70 0 7 FreeSans 80 0 -40 0 GND
port 5 w
flabel metal1 -70 165 -70 165 7 FreeSans 80 0 -40 0 VDD
port 4 w
flabel locali 200 80 200 80 3 FreeSans 80 0 40 0 Y
port 3 e
<< end >>
