magic
tech sky130A
timestamp 1743312914
<< nwell >>
rect -20 45 330 365
<< nmos >>
rect 50 -110 65 -10
rect 115 -110 130 -10
rect 180 -110 195 -10
rect 245 -110 260 -10
<< pmos >>
rect 115 65 130 265
rect 180 65 195 265
<< ndiff >>
rect 0 -25 50 -10
rect 0 -45 15 -25
rect 35 -45 50 -25
rect 0 -75 50 -45
rect 0 -95 15 -75
rect 35 -95 50 -75
rect 0 -110 50 -95
rect 65 -75 115 -10
rect 65 -95 80 -75
rect 100 -95 115 -75
rect 65 -110 115 -95
rect 130 -25 180 -10
rect 130 -45 145 -25
rect 165 -45 180 -25
rect 130 -75 180 -45
rect 130 -95 145 -75
rect 165 -95 180 -75
rect 130 -110 180 -95
rect 195 -25 245 -10
rect 195 -45 210 -25
rect 230 -45 245 -25
rect 195 -110 245 -45
rect 260 -75 310 -10
rect 260 -95 275 -75
rect 295 -95 310 -75
rect 260 -110 310 -95
<< pdiff >>
rect 0 250 115 265
rect 0 230 15 250
rect 35 230 80 250
rect 100 230 115 250
rect 0 200 115 230
rect 0 180 15 200
rect 35 180 80 200
rect 100 180 115 200
rect 0 150 115 180
rect 0 130 15 150
rect 35 130 80 150
rect 100 130 115 150
rect 0 100 115 130
rect 0 80 15 100
rect 35 80 80 100
rect 100 80 115 100
rect 0 65 115 80
rect 130 250 180 265
rect 130 230 145 250
rect 165 230 180 250
rect 130 200 180 230
rect 130 180 145 200
rect 165 180 180 200
rect 130 150 180 180
rect 130 130 145 150
rect 165 130 180 150
rect 130 100 180 130
rect 130 80 145 100
rect 165 80 180 100
rect 130 65 180 80
rect 195 250 310 265
rect 195 230 210 250
rect 230 230 275 250
rect 295 230 310 250
rect 195 200 310 230
rect 195 180 210 200
rect 230 180 275 200
rect 295 180 310 200
rect 195 150 310 180
rect 195 130 210 150
rect 230 130 275 150
rect 295 130 310 150
rect 195 65 310 130
<< ndiffc >>
rect 15 -45 35 -25
rect 15 -95 35 -75
rect 80 -95 100 -75
rect 145 -45 165 -25
rect 145 -95 165 -75
rect 210 -45 230 -25
rect 275 -95 295 -75
<< pdiffc >>
rect 15 230 35 250
rect 80 230 100 250
rect 15 180 35 200
rect 80 180 100 200
rect 15 130 35 150
rect 80 130 100 150
rect 15 80 35 100
rect 80 80 100 100
rect 145 230 165 250
rect 145 180 165 200
rect 145 130 165 150
rect 145 80 165 100
rect 210 230 230 250
rect 275 230 295 250
rect 210 180 230 200
rect 275 180 295 200
rect 210 130 230 150
rect 275 130 295 150
<< psubdiff >>
rect 0 -155 50 -140
rect 0 -175 15 -155
rect 35 -175 50 -155
rect 0 -190 50 -175
rect 130 -155 180 -140
rect 130 -175 145 -155
rect 165 -175 180 -155
rect 130 -190 180 -175
rect 260 -190 310 -140
<< nsubdiff >>
rect 0 295 50 345
rect 130 295 180 345
rect 260 295 310 345
<< psubdiffcont >>
rect 15 -175 35 -155
rect 145 -175 165 -155
<< poly >>
rect 115 265 130 280
rect 180 265 195 280
rect 115 45 130 65
rect 50 35 130 45
rect 50 15 80 35
rect 100 15 130 35
rect 50 5 130 15
rect 50 -10 65 5
rect 115 -10 130 5
rect 180 45 195 65
rect 180 35 260 45
rect 180 15 210 35
rect 230 15 260 35
rect 180 5 260 15
rect 180 -10 195 5
rect 245 -10 260 5
rect 50 -125 65 -110
rect 115 -125 130 -110
rect 180 -125 195 -110
rect 245 -125 260 -110
<< polycont >>
rect 80 15 100 35
rect 210 15 230 35
<< locali >>
rect 5 330 110 340
rect 5 310 15 330
rect 35 310 80 330
rect 100 310 110 330
rect 5 250 110 310
rect 135 330 175 340
rect 135 310 145 330
rect 165 310 175 330
rect 135 300 175 310
rect 200 330 305 340
rect 200 310 210 330
rect 230 310 275 330
rect 295 310 305 330
rect 5 230 15 250
rect 35 230 80 250
rect 100 230 110 250
rect 5 200 110 230
rect 5 180 15 200
rect 35 180 80 200
rect 100 180 110 200
rect 5 150 110 180
rect 5 130 15 150
rect 35 130 80 150
rect 100 130 110 150
rect 5 100 110 130
rect 5 80 15 100
rect 35 80 80 100
rect 100 80 110 100
rect 5 70 110 80
rect 135 250 175 260
rect 135 230 145 250
rect 165 230 175 250
rect 135 200 175 230
rect 135 180 145 200
rect 165 180 175 200
rect 135 150 175 180
rect 135 130 145 150
rect 165 130 175 150
rect 135 100 175 130
rect 200 250 305 310
rect 200 230 210 250
rect 230 230 275 250
rect 295 230 305 250
rect 200 200 305 230
rect 200 180 210 200
rect 230 180 275 200
rect 295 180 305 200
rect 200 150 305 180
rect 200 130 210 150
rect 230 130 275 150
rect 295 130 305 150
rect 200 120 305 130
rect 135 80 145 100
rect 165 90 175 100
rect 165 80 305 90
rect 135 70 305 80
rect 70 35 110 45
rect 70 15 80 35
rect 100 15 110 35
rect 70 5 110 15
rect 200 35 240 45
rect 200 15 210 35
rect 230 15 240 35
rect 200 5 240 15
rect 265 35 305 70
rect 265 15 275 35
rect 295 15 305 35
rect 265 -15 305 15
rect 0 -25 175 -15
rect 0 -45 15 -25
rect 35 -35 145 -25
rect 35 -45 45 -35
rect 0 -75 45 -45
rect 135 -45 145 -35
rect 165 -45 175 -25
rect 0 -95 15 -75
rect 35 -95 45 -75
rect 0 -110 45 -95
rect 70 -75 110 -65
rect 70 -95 80 -75
rect 100 -95 110 -75
rect 5 -155 45 -145
rect 5 -175 15 -155
rect 35 -175 45 -155
rect 5 -185 45 -175
rect 70 -155 110 -95
rect 135 -75 175 -45
rect 200 -25 305 -15
rect 200 -45 210 -25
rect 230 -35 305 -25
rect 230 -45 240 -35
rect 200 -55 240 -45
rect 135 -95 145 -75
rect 165 -85 175 -75
rect 265 -75 305 -65
rect 265 -85 275 -75
rect 165 -95 275 -85
rect 295 -95 305 -75
rect 135 -105 305 -95
rect 70 -175 80 -155
rect 100 -175 110 -155
rect 70 -185 110 -175
rect 135 -155 175 -145
rect 135 -175 145 -155
rect 165 -175 175 -155
rect 135 -185 175 -175
rect 265 -155 305 -145
rect 265 -175 275 -155
rect 295 -175 305 -155
rect 265 -185 305 -175
<< viali >>
rect 15 310 35 330
rect 80 310 100 330
rect 145 310 165 330
rect 210 310 230 330
rect 275 310 295 330
rect 80 15 100 35
rect 210 15 230 35
rect 275 15 295 35
rect 15 -175 35 -155
rect 80 -175 100 -155
rect 145 -175 165 -155
rect 275 -175 295 -155
<< metal1 >>
rect -20 330 330 345
rect -20 310 15 330
rect 35 310 80 330
rect 100 310 145 330
rect 165 310 210 330
rect 230 310 275 330
rect 295 310 330 330
rect -20 295 330 310
rect 70 35 110 45
rect 70 15 80 35
rect 100 15 110 35
rect 70 5 110 15
rect 200 35 240 45
rect 200 15 210 35
rect 230 15 240 35
rect 200 5 240 15
rect 265 35 305 45
rect 265 15 275 35
rect 295 15 305 35
rect 265 5 305 15
rect -20 -155 335 -140
rect -20 -175 15 -155
rect 35 -175 80 -155
rect 100 -175 145 -155
rect 165 -175 275 -155
rect 295 -175 335 -155
rect -20 -190 335 -175
<< labels >>
flabel metal1 70 25 70 25 7 FreeSans 80 0 -40 0 A
port 1 w
flabel metal1 200 25 200 25 7 FreeSans 80 0 -40 0 B
port 2 w
flabel metal1 305 25 305 25 3 FreeSans 80 0 40 0 Y
port 3 e
flabel metal1 -20 320 -20 320 7 FreeSans 80 0 -40 0 VDD
port 4 w
flabel metal1 -20 -165 -20 -165 7 FreeSans 80 0 -40 0 GND
port 5 w
<< end >>
